LIBRARY IEEE ; 
USE IEEE.STD_LOGIC_1164.ALL ; 
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL ; 

entity <your-name> is 
	port(
		); 
end <your-name>;

architecture bhv of <your-name> is 
	component <bla> is
		port(
		);
	end component;

begin

end bhv;

