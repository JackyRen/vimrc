LIBRARY IEEE ; 
USE IEEE.STD_LOGIC_1164.ALL ; 
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL ; 
USE work.GlobalDefines.ALL;

entity <name> is 
	port(
		); 
end <name>;

architecture bhv of <name> is 
	component <bla> is
		port(
		);
	end component;

begin

end bhv;

