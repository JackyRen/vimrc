    component <name> is
        port(

        );
    end component;
